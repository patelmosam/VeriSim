module Not(a, b);
input a;
output b;
assign b = ~a;
endmodule